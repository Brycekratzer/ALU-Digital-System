module storage(

);

endmodule