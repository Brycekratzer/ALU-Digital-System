module adder (
    input [7:0] A,B,
    output reg [7:0]
);
    
endmodule