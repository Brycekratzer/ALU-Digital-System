module operdemux(
    input selector[3:0],
    input val[7:0],
    output reg Y[7:0]
);

// case select or if else statments for each different operation?

endmodule